module curve

import gmp

const (
	zero = gmp.from_u64(0)
	one = gmp.from_u64(1)
	two = gmp.from_u64(2)

	// curve modulo prime for x25519, 2**255 - 19
	cvp_25519 = gmp.from_str('57896044618658097711785492504343953926634992332820282019728792003956564819949')
	// The constant a24 for x25519
	a24_25519 = gmp.from_u64(121665)

	// curve modulo prime for x448 , 2^448 - 2^224 - 1
	cvp_448 = gmp.from_str('726838724295606890549323807888004534353641360687318060281490199180612328166730772686396383698676545930088884461843637361053498018365439') // 2^448 - 2^224 - 1
	// The constant a24 for x448
	a24_448 = gmp.from_u64(39081)

	
)

// y^2 = ax^3 + bx^2 + x mod prime
struct Curve {
	bits_size int
	a24       gmp.Bigint
	prime     gmp.Bigint
}

fn new_x25519_curve() Curve {
	return Curve{
		bits_size: 255
		a24: a24_25519
		prime: cvp_25519
	}
}

fn new_x448_curve() Curve {
	return Curve{
		bits_size: 448
		a24: a24_448
		prime: cvp_448
	}
}

fn new_curve(bits_size int) ?Curve {
	if bits_size !in [255, 448] {
		return error('Bits size $bits_size not permitted, please use 225 or 448')
	}
	mut c := Curve{}
	if bits_size == 255 {
		c = new_x25519_curve()
	}
	if bits_size == 448 {
		c = new_x448_curve()
	}
	return c 
}

fn (cv Curve) x448(mut k []byte, mut u []byte) ?[]byte {
	//first decode k and u and then perform scalar multiply
	//based on formulas from [montgomery].  All calculations are performed modulo p, 
	//and then encode to array of bytes
	if cv.bits_size != 448 && k.len != 56 {
		return error('Bits size should 255 for x25519, but curve has $cv.bits_size')
	}
	_ = k[51]
	mut key := cv.decode_scalar(mut k)?
	mut ucord := cv.decode_x_coordinate(mut u)?

	mut res := cv.scalar_multiply(key, ucord)?
	
	return cv.encode_x_coordinate(mut res)
}

fn (cv Curve) x25519(mut k []byte, mut u []byte) ?[]byte {
	//first decode k and u and then perform scalar multiply
	//based on formulas from [montgomery].  All calculations are performed modulo p, 
	//and then encode to array of bytes
	if cv.bits_size != 255 && k.len != 32 {
		return error('Bits size should 255 for x25519, but curve has $cv.bits_size')
	}
	_ = k[31]
	mut key := cv.decode_scalar(mut k)?
	mut ucord := cv.decode_x_coordinate(mut u)?

	mut res := cv.scalar_multiply(key, ucord)?
	// gmp.clear(mut key)
	// gmp.clear(mut ucord)
	return cv.encode_x_coordinate(mut res)
}

//Scalars are assumed to be randomly generated bytes
fn (cv Curve) decode_scalar(mut k []byte) ?gmp.Bigint {
	if k.len == 0 {
		return error("Not allowed null k length")
	}
	//_ = k[31]
	// mut k := key.clone()
	match cv.bits_size {
		255 {
			//For X25519, in order to decode 32 random bytes as an integer scalar, 
			//set the three least significant bits of the first byte and the most significant bit
   			//of the last to zero, set the second most significant bit of the last
   			//byte to 1 and, finally, decode as little-endian
			_ = k[31]
			k[0] &= 248
			k[31] &= 127
			k[31] |= 64
		}
		448 {
			//for X448, set the two least significant bits of the first byte to 0, and the most
   			//significant bit of the last byte to 1
			_ = k[55]

			k[0] &= 252
			k[55] |= 128
		}
		else {
			return error("k and curve bits size doesn't match")
		}
	}
	return cv.decode_little_endian(k)
}

fn (cv Curve) decode_little_endian(b []byte) ?gmp.Bigint {
	// check if b.len matching with cv.bits
	if b.len !in [32, 56] {
		return error('bytes len $b.len not allowed, please provide valid len bytes')
	}
	match cv.bits_size {
		255 {
			if b.len != 32 {
				return error('bytes len $b.len does not match with underlying curve bits size $cv.bits_size')
			}
		}
		448 {
			if b.len != 56 {
				return error('bytes len $b.len does not match with underlying curve bits size $cv.bits_size')
			}
		}
		else {
			return error('bytes len $b.len does not match with underlying curve bits size $cv.bits_size')
		}
	}
	//_ = b[55]
	mut sum := zero
	for i in 0 .. (cv.bits_size + 7) / 8 {
		mut val := gmp.new()
		// left shift
		gmp.mul_2exp(mut val, gmp.from_u64(b[i]), u64(8 * i))
		sum = sum + val
	}
	return sum
}

fn (cv Curve) decode_x_coordinate(mut u []byte) ?gmp.Bigint {
	//When receiving such an array, implementations of X25519
	//(but not X448) MUST mask the most significant bit in the final byte
	if cv.bits_size % 8 != 0 {
		u[u.len - 1] &= (1 << (cv.bits_size % 8)) - 1
	}
	return cv.decode_little_endian(u)
}

fn (cv Curve) encode_x_coordinate(mut u gmp.Bigint) []byte {
	mut arr := []byte{len: (cv.bits_size + 7) / 8}
	// u = u % cvp_25519
	gmp.mod(mut u, u, cv.prime)

	// placed this allocation out of for loop and call gmp.clear() to release it
	mut val := gmp.new()
	for i in 0 .. arr.len {
		// mut val := gmp.new()
		// this do right shifting
		gmp.tdiv_q_2exp(mut val, u, u64(8 * i))
		// mut d := gmp.new()
		// gmp.and(mut d, val, gmp.from_u64(0xff))
		// arr[i] = byte(d.u64())

		gmp.and(mut val, val, gmp.from_u64(0xff))
		arr[i] = byte(val.u64())
	}
	// gmp.clear(mut val)

	return arr
}

fn (cv Curve) scalar_multiply(k gmp.Bigint, u gmp.Bigint) ?gmp.Bigint {
	if cv.bits_size !in [255, 448] {
		return error("curve bits size doesn't allowed, get $cv.bits_size")
	}
	mut x_1 := u.clone()
	mut x_2 := one
	mut z_2 := zero
	mut x_3 := u.clone()
	mut z_3 := one
	mut swap := zero

	// allocate bigint vars needed for operation outside the loop
	mut k_t := gmp.new()
	mut val := gmp.new()
	mut aa := gmp.new()
	mut bb := gmp.new()
	mut xx := gmp.new()
	for t := cv.bits_size - 1; t >= 0; t-- {
		// this part below, allocated outside for loop
		// mut k_t := gmp.new()
		// mut val := gmp.new()

		// gmp.tdiv_q_2exp(mut val, k, u64(t)) // right shift
		gmp.tdiv_q_2exp(mut val, k, u64(t)) // right shift
		// gmp.and(mut k_t, val, one)
		gmp.and(mut k_t, val, one)
		// mut cs := gmp.new()

		gmp.xor(mut val, swap, k_t)
		// swap = cs
		swap = val

		x_2, x_3 = cswap(swap, x_2, x_3)
		z_2, z_3 = cswap(swap, z_2, z_3)
		swap = k_t

		mut a := (x_2 + z_2) % cv.prime
		// mut aa := gmp.new()
		// eliminate a allocation
		gmp.powm_sec(mut aa, a, curve.two, cv.prime)

		mut b := (x_2 - z_2) % cv.prime
		// mut bb := gmp.new()
		gmp.powm_sec(mut bb, b, curve.two, cv.prime)

		mut e := (aa - bb) % cv.prime
		mut c := (x_3 + z_3) % cv.prime
		mut d := (x_3 - z_3) % cv.prime

		mut da := (d * a) % cv.prime
		mut cb := (c * b) % cv.prime

		gmp.powm_sec(mut x_3, (da + cb) % cv.prime, curve.two, cv.prime)
		// mut xx := gmp.new()
		gmp.powm_sec(mut xx, (da - cb) % cv.prime, curve.two, cv.prime)

		// z_3 = (x_1 * xx) % cv.prime
		z_3 = (x_1 * xx) % cv.prime
		x_2 = (aa * bb) % cv.prime
		z_2 = e * ((aa + (cv.a24 * e) % cv.prime) % cv.prime)
	}
	x_2, x_3 = cswap(swap, x_2, x_3)
	z_2, z_3 = cswap(swap, z_2, z_3)
	// mut zz := gmp.new()
	// gmp.powm(mut zz, z_2, cv.prime - two, cv.prime)
	gmp.powm_sec(mut val, z_2, cv.prime - curve.two, cv.prime)

	// res := (x_2 * zz) % cv.prime
	res := (x_2 * val) % cv.prime

	return res
}

fn cswap(swap gmp.Bigint, x_2 gmp.Bigint, x_3 gmp.Bigint) (gmp.Bigint, gmp.Bigint) {
	mask := zero - swap
	mut dummy := gmp.new()
	mut vv := gmp.new()
	gmp.xor(mut vv, x_2, x_3)
	gmp.and(mut dummy, mask, vv)
	mut r1 := gmp.new()
	mut r2 := gmp.new()

	gmp.xor(mut r1, x_2, dummy)
	gmp.xor(mut r2, x_3, dummy)

	return r1, r2
}
